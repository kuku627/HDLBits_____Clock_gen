module top_module(
    input a,b,
    output sum,cout
);
assign cout=a&b;
assign sum=a^b;


endmodule