module top_module (
    input a,
    input b,
    output wire q );
    


assign q=a&b;

endmodule